// board_kernel_interface.v

// Generated using ACDS version 19.1 240

`timescale 1 ps / 1 ps
module board_kernel_interface (
		input  wire        kernel_cra_waitrequest,        //               kernel_cra.waitrequest
		input  wire [63:0] kernel_cra_readdata,           //                         .readdata
		input  wire        kernel_cra_readdatavalid,      //                         .readdatavalid
		output wire [0:0]  kernel_cra_burstcount,         //                         .burstcount
		output wire [63:0] kernel_cra_writedata,          //                         .writedata
		output wire [29:0] kernel_cra_address,            //                         .address
		output wire        kernel_cra_write,              //                         .write
		output wire        kernel_cra_read,               //                         .read
		output wire [7:0]  kernel_cra_byteenable,         //                         .byteenable
		output wire        kernel_cra_debugaccess,        //                         .debugaccess
		output wire        ctrl_waitrequest,              //                     ctrl.waitrequest
		output wire [31:0] ctrl_readdata,                 //                         .readdata
		output wire        ctrl_readdatavalid,            //                         .readdatavalid
		input  wire [0:0]  ctrl_burstcount,               //                         .burstcount
		input  wire [31:0] ctrl_writedata,                //                         .writedata
		input  wire [13:0] ctrl_address,                  //                         .address
		input  wire        ctrl_write,                    //                         .write
		input  wire        ctrl_read,                     //                         .read
		input  wire [3:0]  ctrl_byteenable,               //                         .byteenable
		input  wire        ctrl_debugaccess,              //                         .debugaccess
		output wire [1:0]  acl_bsp_memorg_host0x018_mode, // acl_bsp_memorg_host0x018.mode
		input  wire        clk_clk,                       //                      clk.clk
		input  wire        reset_reset_n,                 //                    reset.reset_n
		input  wire [0:0]  kernel_irq_from_kernel_irq,    //   kernel_irq_from_kernel.irq
		output wire        kernel_irq_to_host_irq,        //       kernel_irq_to_host.irq
		input  wire        sw_reset_in_reset,             //              sw_reset_in.reset
		input  wire        kernel_clk_clk,                //               kernel_clk.clk
		output wire        kernel_reset_reset_n,          //             kernel_reset.reset_n
		output wire        sw_reset_export_reset_n        //          sw_reset_export.reset_n
	);

	board_kernel_interface_kernel_interface_151_5tpfcyy kernel_interface (
		.kernel_cra_waitrequest        (kernel_cra_waitrequest),        //   input,   width = 1,               kernel_cra.waitrequest
		.kernel_cra_readdata           (kernel_cra_readdata),           //   input,  width = 64,                         .readdata
		.kernel_cra_readdatavalid      (kernel_cra_readdatavalid),      //   input,   width = 1,                         .readdatavalid
		.kernel_cra_burstcount         (kernel_cra_burstcount),         //  output,   width = 1,                         .burstcount
		.kernel_cra_writedata          (kernel_cra_writedata),          //  output,  width = 64,                         .writedata
		.kernel_cra_address            (kernel_cra_address),            //  output,  width = 30,                         .address
		.kernel_cra_write              (kernel_cra_write),              //  output,   width = 1,                         .write
		.kernel_cra_read               (kernel_cra_read),               //  output,   width = 1,                         .read
		.kernel_cra_byteenable         (kernel_cra_byteenable),         //  output,   width = 8,                         .byteenable
		.kernel_cra_debugaccess        (kernel_cra_debugaccess),        //  output,   width = 1,                         .debugaccess
		.ctrl_waitrequest              (ctrl_waitrequest),              //  output,   width = 1,                     ctrl.waitrequest
		.ctrl_readdata                 (ctrl_readdata),                 //  output,  width = 32,                         .readdata
		.ctrl_readdatavalid            (ctrl_readdatavalid),            //  output,   width = 1,                         .readdatavalid
		.ctrl_burstcount               (ctrl_burstcount),               //   input,   width = 1,                         .burstcount
		.ctrl_writedata                (ctrl_writedata),                //   input,  width = 32,                         .writedata
		.ctrl_address                  (ctrl_address),                  //   input,  width = 14,                         .address
		.ctrl_write                    (ctrl_write),                    //   input,   width = 1,                         .write
		.ctrl_read                     (ctrl_read),                     //   input,   width = 1,                         .read
		.ctrl_byteenable               (ctrl_byteenable),               //   input,   width = 4,                         .byteenable
		.ctrl_debugaccess              (ctrl_debugaccess),              //   input,   width = 1,                         .debugaccess
		.acl_bsp_memorg_host0x018_mode (acl_bsp_memorg_host0x018_mode), //  output,   width = 2, acl_bsp_memorg_host0x018.mode
		.clk_clk                       (clk_clk),                       //   input,   width = 1,                      clk.clk
		.reset_reset_n                 (reset_reset_n),                 //   input,   width = 1,                    reset.reset_n
		.kernel_irq_from_kernel_irq    (kernel_irq_from_kernel_irq),    //   input,   width = 1,   kernel_irq_from_kernel.irq
		.kernel_irq_to_host_irq        (kernel_irq_to_host_irq),        //  output,   width = 1,       kernel_irq_to_host.irq
		.sw_reset_in_reset             (sw_reset_in_reset),             //   input,   width = 1,              sw_reset_in.reset
		.kernel_clk_clk                (kernel_clk_clk),                //   input,   width = 1,               kernel_clk.clk
		.kernel_reset_reset_n          (kernel_reset_reset_n),          //  output,   width = 1,             kernel_reset.reset_n
		.sw_reset_export_reset_n       (sw_reset_export_reset_n)        //  output,   width = 1,          sw_reset_export.reset_n
	);

endmodule
